`timescale 1ns/1ps

module tb_instruction_decode();

endmodule