module PC_MUX_ENUM();
    localparam [1:0] NOP = 2'b00;
    localparam [1:0] PC_ADDER = 2'b01;
    localparam [1:0] ALU_OUT = 2'b10;
endmodule