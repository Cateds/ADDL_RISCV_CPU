module reg_if_id(
        // * Clock Sync Signals Connection --------------------
        input clk,
        input rst_n,
        // * Pipeline Signals Connection --------------------
        input stall,
        input flush,
        // * Input Signals Connection --------------------

        // * Output Signals Connection --------------------
    );
endmodule
