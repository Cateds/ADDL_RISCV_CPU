module memory_operation();
endmodule