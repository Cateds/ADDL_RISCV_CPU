module PC_MUX_ENUM();
    parameter NOP = 2'b00;
    parameter PC_ADDER = 2'b01;
    parameter ALU_OUT = 2'b10;
endmodule