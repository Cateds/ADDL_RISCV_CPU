module execute();
endmodule