module instruction_fetch(
        // * Clock Sync Signals Connection --------------------
        input wire clk,
        input wire rst_n,

        // * Internal Signals Connection --------------------
        input wire [1:0] branch,
        input wire [31:0] alu_result,
        input wire [31:0] pc_adder_result,

        output wire [31:0] pc,
        output wire [31:0] pc_next,
        output wire [31:0] instruction,

        // * External Signals Connection --------------------
        output wire [31:0] rom_addr,
        input wire [31:0] rom_data,
        output wire rom_en
    );

    // output declaration of module program_counter
    program_counter
        u_program_counter(
            .branch          	(branch           ),
            .en              	(en               ),
            .clk             	(clk              ),
            .rst_n           	(rst_n            ),
            .alu_result      	(alu_result       ),
            .pc_adder_result 	(pc_adder_result  ),
            .pc              	(pc               ),
            .pc_next         	(pc_next          )
        );

    assign rom_addr = pc; // PC作为ROM的地址
    assign instruction = rom_data; // 从ROM中读取指令
    assign rom_en = 1'b1;
endmodule
