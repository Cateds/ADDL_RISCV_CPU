module gpio(
    // ----- Clock Sync Signals Connection -----
    input wire clk,
    input wire rst_n,
    input wire gpio_ce,

    // ----- Internal Signals Connection -----
    input wire bus_we,
    input wire bus_re,
    

    // ----- External Signals Connection -----
);
endmodule